library



entity SignExtend is
port(x:in std_logic_vector(15 downto 0);y:out std_logic_vector(31 downto 0));
end SignExtend;

